module ArrayMultiplier4 (
    input [3:0] A,
    input [3:0] B,
    output [7:0] Prod
);

    // Generate Product using nested loops
    generate
        for (genvar i = 0; i < 4; i = i + 1) begin : gen_mult
            for (genvar j = 0; j < 4; j = j + 1) begin : gen_add
                assign Prod[i + j] = A[i] & B[j];
            end
        end
    endgenerate

endmodule
